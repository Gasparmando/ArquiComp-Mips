`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:29:01 02/02/2020 
// Design Name: 
// Module Name:    MEM_MemoryAccess 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module _4_MEM_MemoryAccess(
    );

DataMemory dm();

MEM_WB mem_wb();

endmodule
